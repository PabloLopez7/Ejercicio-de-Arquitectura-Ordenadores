----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:41:03 05/23/2022 
-- Design Name: 
-- Module Name:    Promedio1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Promedio1 is
    Port ( A,B : in  STD_LOGIC (0 downto 3);
           C : out  STD_LOGIC(0 downto 3));
end Promedio1;

architecture Behavioral of Promedio1 is

begin


end Behavioral;

