----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:46:04 05/23/2022 
-- Design Name: 
-- Module Name:    MUX - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity MUX is
    Port ( E0,E1,E2,E3 : in  STD_LOGIC;
           S0,S1 : in  STD_LOGIC;
           F : out  STD_LOGIC);
end MUX;

architecture Behavioral of MUX is

begin


end Behavioral;

