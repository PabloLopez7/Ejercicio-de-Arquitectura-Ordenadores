----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:33:53 05/23/2022 
-- Design Name: 
-- Module Name:    Proyecto - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Proyecto is
    Port ( P0 : in      STD_LOGIC;
           P1 : in      STD_LOGIC;
           P2 : in      STD_LOGIC;
           X :  buffer  STD_LOGIC;
           A1 : out     STD_LOGIC;
           A2 : out     STD_LOGIC);
end Proyecto;

architecture Behavioral of Proyecto is

begin


end Behavioral;

