----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:13:38 05/23/2022 
-- Design Name: 
-- Module Name:    ejemplos - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ejemplos is
    Port ( x1 : in  STD_LOGIC;
           x2 : in  STD_LOGIC;
           fa : out  STD_LOGIC;
           fb : out  STD_LOGIC);
end ejemplos;

architecture Behavioral of ejemplos is

begin


end Behavioral;

